--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   13:32:59 06/16/2015
-- Design Name:   
-- Module Name:   C:/project10/MUX_tb.vhd
-- Project Name:  project10
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: MUX
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY MUX_tb IS
END MUX_tb;
 
ARCHITECTURE behavior OF MUX_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT MUX
    PORT(
         mode : IN  std_logic;
         next_add : IN  std_logic_vector(4 downto 0);
         op_addr : IN  std_logic_vector(4 downto 0);
         out_add : OUT  std_logic_vector(4 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal mode : std_logic := '0';
   signal next_add : std_logic_vector(4 downto 0) := (others => '0');
   signal op_addr : std_logic_vector(4 downto 0) := (others => '0');

 	--Outputs
   signal out_add : std_logic_vector(4 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: MUX PORT MAP (
          mode => mode,
          next_add => next_add,
          op_addr => op_addr,
          out_add => out_add
        );

 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 20 ns;	
			mode<='0';
			next_add<="00010";
			op_addr<="01010";
		wait for 20 ns;	
			mode<='1';
			next_add<="00010";
			op_addr<="01010";
		wait for 20 ns;	
			next_add<="00011";
			op_addr<="01000";
		wait for 20 ns;	
			mode<='0';
			next_add<="00011";
			op_addr<="01000";

      -- insert stimulus here 

      wait;
   end process;

END;
